module submodule03 (
  // Clock and reset
  input  wire  clk,
  input  wire                rst_n
);


endmodule